module dcdw23_module (
    
);
    input clk, rst;
    input [15:0]

endmodule //dcdw23_module